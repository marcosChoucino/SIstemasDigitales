library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity LCD_DRAWING IS
	port
	(	--entradas
		reset,CLK		: in std_logic;
		DEL_SCREEN, DRAW_FIG	: in std_logic;
		COLOUR_CODE		: in std_logic_vector(2 downto 0);
		DONE_CURSOR,DONE_COLOUR	: in std_logic;

		--salidas
		OP_SETCURSOR		: out std_logic;
		XCOL			: out std_logic_vector(7 downto 0);
		YROW			: out std_logic_vector(8 downto 0);
		OP_DRAWCOLOUR	: out std_logic;
		RGB			: out std_logic_vector(15 downto 0);
		NUMPIX			: out std_logic_vector(16 downto 0)
	);
end LCD_DRAWING;


architecture ARCH_LCD_DRAWING of LCD_DRAWING is

	type state is (E0,E1,E2,E3,E4,E5,E6,E7,E8);
	signal EP,ES: state;

	--se�ales registro colores
	signal COLOUR_CODE_OUT : unsigned(2 downto 0);
	signal LD_COLOUR		: std_logic;
	--contador colorines
	signal TC_DIAG	:  	std_logic;
	signal OUT_DIAG :	unsigned(7 downto 0);
	signal LD_DIAG : 	std_logic;
	signal INC_DIAG : 	std_logic;
	--contador YROW
	signal YROW2	:  	unsigned(8 downto 0);
	signal LD_Y : 	std_logic;
	signal INC_Y : 	std_logic;
	--contador XCOL
	signal XCOL2	:  	unsigned(7 downto 0);
	signal LD_X : 	std_logic;
	signal INC_X : 	std_logic;
	--contador numpix

	signal BORRAR_DIAGONAL: std_logic;

begin
-------------------------------------------------------------------------------------------
	-- CONTROL UNIT
-------------------------------------------------------------------------------------------
	--
	-- Current state Register (State Machine)
	process (CLK, reset)
	begin
		if reset = '1' then EP <= E0;
	  	elsif rising_edge(CLK) then EP <= ES ;
		end if;
	end process;

	-- Next state generation logic
	process (EP,DEL_SCREEN,DRAW_FIG,DONE_CURSOR,DONE_COLOUR,TC_DIAG)
	begin
  		case EP is
			when E0 => 	if (DEL_SCREEN='0' and DRAW_FIG='0') then ES <= E0;          	-- |
	           			elsif (DEL_SCREEN='1') then ES <= E1;         			-- |Initial state
                   	elsif (DRAW_FIG='1') then ES <= E4; 				-- |
							else ES <= E0;                                   		-- |
	       	   			end if;
			--DEL_SCREEN
			when E1 => ES <= E2;       
			when E2 => 	if(DONE_CURSOR='1')then ES <= E3;
					else ES <= E2; --handsake done_cursor_delScreen
					end if;
					         
			when E3 => 	if(DONE_COLOUR='1')then ES <= E0;
					else ES <= E3; --handsake done_colour_delScreen 
					end if;
                  	--DRAW_FIG
			when E4 => ES <= E5;                                                    
			when E5 => ES <= E6;                         
			when E6 =>	if(DONE_CURSOR='1')then ES <= E7;
					else ES <= E5; --handsake done_cursor_DRAW_FIG
					end if;
			when E7 => 	if(DONE_COLOUR='1' and TC_DIAG='1')then ES <= E0;
					elsif(DONE_COLOUR='1' and TC_DIAG='0')then ES <= E8; --handsake done_colour_DRAW_FIG
					else ES <= E7;  
					end if;     
			when E8 => ES <= E5;
  		end case;
	end process;
	
	-- Control signals generation logic
	LD_X <= '1' when (EP=E1 or EP=E4) else '0';
	LD_Y <= '1' when (EP=E1 or EP=E4) else '0';
	LD_COLOUR <= '1' when (EP=E1 or EP=E4) else '0';
	LD_DIAG <= '1' when (EP=E4) else '0';
	OP_DRAWCOLOUR <= '1' when(EP=E3 or EP=E7) else '0';
	OP_SETCURSOR <= '1' when(EP=E2 or EP=E6) else '0';	
	BORRAR_DIAGONAL <= '1' when (EP=E2 or EP=E1) else '0'; -- tal vez mejor en E1 o en los dos
	INC_DIAG <= '1' when (EP=E5) else '0';
	INC_Y<= '1' when (EP=E8) else '0';
	INC_X<= '1' when (EP=E8) else '0';

-------------------------------------------------------------------------------------------
-- PROCESS UNIT
-------------------------------------------------------------------------------------------
	
--------------------------------------------
--REGISTRO COLORES
--------------------------------------------
	--registro que seleccionara los colores 
	process(CLK,reset)
	begin
	if (reset='1') then COLOUR_CODE_OUT <=(others=>'0');
   	elsif rising_edge(CLK) then 
	     	if (LD_COLOUR='1') then COLOUR_CODE_OUT <= unsigned(COLOUR_CODE);
         end if;
	end if;		  
	end process;
	
--------------------------------------------
--REGISTRO CONTADOR DIAGONAL
--------------------------------------------
	process(CLK,reset)
	begin
		if (reset='1') then OUT_DIAG<= x"F0"; TC_DIAG<='0'; 
   	elsif rising_edge(CLK) then 
           	if (INC_DIAG='1') then OUT_DIAG <= OUT_DIAG - 1;
            elsif (LD_DIAG ='1') then OUT_DIAG <= x"F0";
            end if;
				if(OUT_DIAG=x"00") then TC_DIAG<='1';
				else TC_DIAG<='0';
				end if;
		end if;		  
	end process;

--------------------------------------------
--REGISTRO CONTADOR YROW
--------------------------------------------
	process(CLK,reset)
	begin
		if (reset='1') then YROW2<=(others=>'0');
   		elsif rising_edge(CLK) then 
	   		if (INC_Y='1') then YROW2 <= YROW2 + 1;
            		elsif (LD_Y ='1') then YROW2 <= "000000000";
            		end if;
		end if;		  
	end process;
	YROW <=std_logic_vector(YROW2);
--------------------------------------------
--REGISTRO CONTADOR XCOL
--------------------------------------------
	process(CLK,reset)
	begin
		if (reset='1') then XCOL2<=(others=>'0');
   		elsif rising_edge(CLK) then 
	   		if (INC_X='1') then XCOL2 <= XCOL2 + 1;
            		elsif (LD_X ='1') then XCOL2 <= "00000000";
            		end if;
		end if;		  
	end process;
	XCOL <= std_logic_vector(XCOL2);
--------------------------------------------
--MULTIFLEXOR DE LOS COLORES :p
--------------------------------------------
 
-- RGB 8:1 Multiplexer
	RGB <= x"F81F" when COLOUR_CODE_OUT="000" else    -- ROJO 
	 		x"001F" when COLOUR_CODE_OUT="001" else   -- AZUL
           			x"07E0" when COLOUR_CODE_OUT="010" else   -- VERDE
			x"FFE0" when COLOUR_CODE_OUT="011" else	-- AMARILLO
           	 		x"F81F" when COLOUR_CODE_OUT="100" else -- ROSA
            		x"07FF" when COLOUR_CODE_OUT="101" else    -- CYAN
            		x"FFFF" when COLOUR_CODE_OUT="110" else   --BLANCO
            		x"0000";		-- NEGRO



--------------------------------------------
--MULTIFLEXOR NUMPIX
--------------------------------------------

NUMPIX <= "00000000000000001" when BORRAR_DIAGONAL = '0' else "10010110000000000";
end ARCH_LCD_DRAWING;						


	